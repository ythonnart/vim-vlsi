--------------------------------------------------------------------------------
-- Compilation test
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Scratchpad, don't remove marker
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
-- begin scratchpad

-- end scratchpad
